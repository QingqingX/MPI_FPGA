// nios2.v

// Generated using ACDS version 15.1 185

`timescale 1 ps / 1 ps
module nios2 (
		output wire [127:0] acc_0_packet_out_packet,   //   acc_0_packet_out.packet
		output wire         acc_0_packet_out_valid,    //                   .valid
		input  wire [127:0] acc_recv_0_pack_in_packet, // acc_recv_0_pack_in.packet
		input  wire         acc_recv_0_pack_in_valid,  //                   .valid
		input  wire         clk_clk,                   //                clk.clk
		input  wire         reset_reset_n              //              reset.reset_n
	);

	wire         pll_0_outclk0_clk;                                                          // pll_0:outclk_0 -> [arbit_0:clk, irq_mapper:clk, jtaguart_0:clk, mem:clk, mem:clk2, mm_interconnect_0:pll_0_outclk0_clk, mm_interconnect_1:pll_0_outclk0_clk, nios2_0:clk, performance_counter_0:clk, rst_controller:clk, sys_clk_timer:clk, sysid:clock]
	wire  [31:0] acc_recv_0_conduit_end_write_addr;                                          // acc_recv_0:write_addr -> arbit_0:write_addr_r
	wire         acc_recv_0_conduit_end_write;                                               // acc_recv_0:write -> arbit_0:write_r
	wire  [31:0] acc_recv_0_conduit_end_data_to_mem;                                         // acc_recv_0:data_to_mem -> arbit_0:data_to_mem_r
	wire  [31:0] nios2_0_custom_instruction_master_multi_dataa;                              // nios2_0:A_ci_multi_dataa -> nios2_0_custom_instruction_master_translator:ci_slave_multi_dataa
	wire         nios2_0_custom_instruction_master_multi_writerc;                            // nios2_0:A_ci_multi_writerc -> nios2_0_custom_instruction_master_translator:ci_slave_multi_writerc
	wire  [31:0] nios2_0_custom_instruction_master_multi_result;                             // nios2_0_custom_instruction_master_translator:ci_slave_multi_result -> nios2_0:A_ci_multi_result
	wire         nios2_0_custom_instruction_master_clk;                                      // nios2_0:A_ci_multi_clock -> nios2_0_custom_instruction_master_translator:ci_slave_multi_clk
	wire  [31:0] nios2_0_custom_instruction_master_multi_datab;                              // nios2_0:A_ci_multi_datab -> nios2_0_custom_instruction_master_translator:ci_slave_multi_datab
	wire         nios2_0_custom_instruction_master_start;                                    // nios2_0:A_ci_multi_start -> nios2_0_custom_instruction_master_translator:ci_slave_multi_start
	wire   [4:0] nios2_0_custom_instruction_master_multi_b;                                  // nios2_0:A_ci_multi_b -> nios2_0_custom_instruction_master_translator:ci_slave_multi_b
	wire   [4:0] nios2_0_custom_instruction_master_multi_c;                                  // nios2_0:A_ci_multi_c -> nios2_0_custom_instruction_master_translator:ci_slave_multi_c
	wire         nios2_0_custom_instruction_master_reset_req;                                // nios2_0:A_ci_multi_reset_req -> nios2_0_custom_instruction_master_translator:ci_slave_multi_reset_req
	wire         nios2_0_custom_instruction_master_done;                                     // nios2_0_custom_instruction_master_translator:ci_slave_multi_done -> nios2_0:A_ci_multi_done
	wire   [4:0] nios2_0_custom_instruction_master_multi_a;                                  // nios2_0:A_ci_multi_a -> nios2_0_custom_instruction_master_translator:ci_slave_multi_a
	wire         nios2_0_custom_instruction_master_clk_en;                                   // nios2_0:A_ci_multi_clk_en -> nios2_0_custom_instruction_master_translator:ci_slave_multi_clken
	wire         nios2_0_custom_instruction_master_reset;                                    // nios2_0:A_ci_multi_reset -> nios2_0_custom_instruction_master_translator:ci_slave_multi_reset
	wire         nios2_0_custom_instruction_master_multi_readrb;                             // nios2_0:A_ci_multi_readrb -> nios2_0_custom_instruction_master_translator:ci_slave_multi_readrb
	wire         nios2_0_custom_instruction_master_multi_readra;                             // nios2_0:A_ci_multi_readra -> nios2_0_custom_instruction_master_translator:ci_slave_multi_readra
	wire   [7:0] nios2_0_custom_instruction_master_multi_n;                                  // nios2_0:A_ci_multi_n -> nios2_0_custom_instruction_master_translator:ci_slave_multi_n
	wire         nios2_0_custom_instruction_master_translator_multi_ci_master_readra;        // nios2_0_custom_instruction_master_translator:multi_ci_master_readra -> nios2_0_custom_instruction_master_multi_xconnect:ci_slave_readra
	wire   [4:0] nios2_0_custom_instruction_master_translator_multi_ci_master_a;             // nios2_0_custom_instruction_master_translator:multi_ci_master_a -> nios2_0_custom_instruction_master_multi_xconnect:ci_slave_a
	wire   [4:0] nios2_0_custom_instruction_master_translator_multi_ci_master_b;             // nios2_0_custom_instruction_master_translator:multi_ci_master_b -> nios2_0_custom_instruction_master_multi_xconnect:ci_slave_b
	wire         nios2_0_custom_instruction_master_translator_multi_ci_master_clk;           // nios2_0_custom_instruction_master_translator:multi_ci_master_clk -> nios2_0_custom_instruction_master_multi_xconnect:ci_slave_clk
	wire         nios2_0_custom_instruction_master_translator_multi_ci_master_readrb;        // nios2_0_custom_instruction_master_translator:multi_ci_master_readrb -> nios2_0_custom_instruction_master_multi_xconnect:ci_slave_readrb
	wire   [4:0] nios2_0_custom_instruction_master_translator_multi_ci_master_c;             // nios2_0_custom_instruction_master_translator:multi_ci_master_c -> nios2_0_custom_instruction_master_multi_xconnect:ci_slave_c
	wire         nios2_0_custom_instruction_master_translator_multi_ci_master_start;         // nios2_0_custom_instruction_master_translator:multi_ci_master_start -> nios2_0_custom_instruction_master_multi_xconnect:ci_slave_start
	wire         nios2_0_custom_instruction_master_translator_multi_ci_master_reset_req;     // nios2_0_custom_instruction_master_translator:multi_ci_master_reset_req -> nios2_0_custom_instruction_master_multi_xconnect:ci_slave_reset_req
	wire         nios2_0_custom_instruction_master_translator_multi_ci_master_done;          // nios2_0_custom_instruction_master_multi_xconnect:ci_slave_done -> nios2_0_custom_instruction_master_translator:multi_ci_master_done
	wire   [7:0] nios2_0_custom_instruction_master_translator_multi_ci_master_n;             // nios2_0_custom_instruction_master_translator:multi_ci_master_n -> nios2_0_custom_instruction_master_multi_xconnect:ci_slave_n
	wire  [31:0] nios2_0_custom_instruction_master_translator_multi_ci_master_result;        // nios2_0_custom_instruction_master_multi_xconnect:ci_slave_result -> nios2_0_custom_instruction_master_translator:multi_ci_master_result
	wire         nios2_0_custom_instruction_master_translator_multi_ci_master_clk_en;        // nios2_0_custom_instruction_master_translator:multi_ci_master_clken -> nios2_0_custom_instruction_master_multi_xconnect:ci_slave_clken
	wire  [31:0] nios2_0_custom_instruction_master_translator_multi_ci_master_datab;         // nios2_0_custom_instruction_master_translator:multi_ci_master_datab -> nios2_0_custom_instruction_master_multi_xconnect:ci_slave_datab
	wire  [31:0] nios2_0_custom_instruction_master_translator_multi_ci_master_dataa;         // nios2_0_custom_instruction_master_translator:multi_ci_master_dataa -> nios2_0_custom_instruction_master_multi_xconnect:ci_slave_dataa
	wire         nios2_0_custom_instruction_master_translator_multi_ci_master_reset;         // nios2_0_custom_instruction_master_translator:multi_ci_master_reset -> nios2_0_custom_instruction_master_multi_xconnect:ci_slave_reset
	wire         nios2_0_custom_instruction_master_translator_multi_ci_master_writerc;       // nios2_0_custom_instruction_master_translator:multi_ci_master_writerc -> nios2_0_custom_instruction_master_multi_xconnect:ci_slave_writerc
	wire         nios2_0_custom_instruction_master_multi_xconnect_ci_master0_readra;         // nios2_0_custom_instruction_master_multi_xconnect:ci_master0_readra -> nios2_0_custom_instruction_master_multi_slave_translator0:ci_slave_readra
	wire   [4:0] nios2_0_custom_instruction_master_multi_xconnect_ci_master0_a;              // nios2_0_custom_instruction_master_multi_xconnect:ci_master0_a -> nios2_0_custom_instruction_master_multi_slave_translator0:ci_slave_a
	wire   [4:0] nios2_0_custom_instruction_master_multi_xconnect_ci_master0_b;              // nios2_0_custom_instruction_master_multi_xconnect:ci_master0_b -> nios2_0_custom_instruction_master_multi_slave_translator0:ci_slave_b
	wire         nios2_0_custom_instruction_master_multi_xconnect_ci_master0_readrb;         // nios2_0_custom_instruction_master_multi_xconnect:ci_master0_readrb -> nios2_0_custom_instruction_master_multi_slave_translator0:ci_slave_readrb
	wire   [4:0] nios2_0_custom_instruction_master_multi_xconnect_ci_master0_c;              // nios2_0_custom_instruction_master_multi_xconnect:ci_master0_c -> nios2_0_custom_instruction_master_multi_slave_translator0:ci_slave_c
	wire         nios2_0_custom_instruction_master_multi_xconnect_ci_master0_clk;            // nios2_0_custom_instruction_master_multi_xconnect:ci_master0_clk -> nios2_0_custom_instruction_master_multi_slave_translator0:ci_slave_clk
	wire  [31:0] nios2_0_custom_instruction_master_multi_xconnect_ci_master0_ipending;       // nios2_0_custom_instruction_master_multi_xconnect:ci_master0_ipending -> nios2_0_custom_instruction_master_multi_slave_translator0:ci_slave_ipending
	wire         nios2_0_custom_instruction_master_multi_xconnect_ci_master0_start;          // nios2_0_custom_instruction_master_multi_xconnect:ci_master0_start -> nios2_0_custom_instruction_master_multi_slave_translator0:ci_slave_start
	wire         nios2_0_custom_instruction_master_multi_xconnect_ci_master0_reset_req;      // nios2_0_custom_instruction_master_multi_xconnect:ci_master0_reset_req -> nios2_0_custom_instruction_master_multi_slave_translator0:ci_slave_reset_req
	wire         nios2_0_custom_instruction_master_multi_xconnect_ci_master0_done;           // nios2_0_custom_instruction_master_multi_slave_translator0:ci_slave_done -> nios2_0_custom_instruction_master_multi_xconnect:ci_master0_done
	wire   [7:0] nios2_0_custom_instruction_master_multi_xconnect_ci_master0_n;              // nios2_0_custom_instruction_master_multi_xconnect:ci_master0_n -> nios2_0_custom_instruction_master_multi_slave_translator0:ci_slave_n
	wire  [31:0] nios2_0_custom_instruction_master_multi_xconnect_ci_master0_result;         // nios2_0_custom_instruction_master_multi_slave_translator0:ci_slave_result -> nios2_0_custom_instruction_master_multi_xconnect:ci_master0_result
	wire         nios2_0_custom_instruction_master_multi_xconnect_ci_master0_estatus;        // nios2_0_custom_instruction_master_multi_xconnect:ci_master0_estatus -> nios2_0_custom_instruction_master_multi_slave_translator0:ci_slave_estatus
	wire         nios2_0_custom_instruction_master_multi_xconnect_ci_master0_clk_en;         // nios2_0_custom_instruction_master_multi_xconnect:ci_master0_clken -> nios2_0_custom_instruction_master_multi_slave_translator0:ci_slave_clken
	wire  [31:0] nios2_0_custom_instruction_master_multi_xconnect_ci_master0_datab;          // nios2_0_custom_instruction_master_multi_xconnect:ci_master0_datab -> nios2_0_custom_instruction_master_multi_slave_translator0:ci_slave_datab
	wire  [31:0] nios2_0_custom_instruction_master_multi_xconnect_ci_master0_dataa;          // nios2_0_custom_instruction_master_multi_xconnect:ci_master0_dataa -> nios2_0_custom_instruction_master_multi_slave_translator0:ci_slave_dataa
	wire         nios2_0_custom_instruction_master_multi_xconnect_ci_master0_reset;          // nios2_0_custom_instruction_master_multi_xconnect:ci_master0_reset -> nios2_0_custom_instruction_master_multi_slave_translator0:ci_slave_reset
	wire         nios2_0_custom_instruction_master_multi_xconnect_ci_master0_writerc;        // nios2_0_custom_instruction_master_multi_xconnect:ci_master0_writerc -> nios2_0_custom_instruction_master_multi_slave_translator0:ci_slave_writerc
	wire  [31:0] nios2_0_custom_instruction_master_multi_slave_translator0_ci_master_result; // acc_0:result -> nios2_0_custom_instruction_master_multi_slave_translator0:ci_master_result
	wire         nios2_0_custom_instruction_master_multi_slave_translator0_ci_master_clk;    // nios2_0_custom_instruction_master_multi_slave_translator0:ci_master_clk -> acc_0:nios_clk
	wire         nios2_0_custom_instruction_master_multi_slave_translator0_ci_master_clk_en; // nios2_0_custom_instruction_master_multi_slave_translator0:ci_master_clken -> acc_0:clk_en
	wire  [31:0] nios2_0_custom_instruction_master_multi_slave_translator0_ci_master_datab;  // nios2_0_custom_instruction_master_multi_slave_translator0:ci_master_datab -> acc_0:data_in_b
	wire  [31:0] nios2_0_custom_instruction_master_multi_slave_translator0_ci_master_dataa;  // nios2_0_custom_instruction_master_multi_slave_translator0:ci_master_dataa -> acc_0:data_in_a
	wire         nios2_0_custom_instruction_master_multi_slave_translator0_ci_master_start;  // nios2_0_custom_instruction_master_multi_slave_translator0:ci_master_start -> acc_0:start
	wire         nios2_0_custom_instruction_master_multi_slave_translator0_ci_master_reset;  // nios2_0_custom_instruction_master_multi_slave_translator0:ci_master_reset -> acc_0:reset
	wire         nios2_0_custom_instruction_master_multi_slave_translator0_ci_master_done;   // acc_0:done -> nios2_0_custom_instruction_master_multi_slave_translator0:ci_master_done
	wire   [2:0] nios2_0_custom_instruction_master_multi_slave_translator0_ci_master_n;      // nios2_0_custom_instruction_master_multi_slave_translator0:ci_master_n -> acc_0:in_opcode
	wire         nios2_0_custom_instruction_master_multi_xconnect_ci_master1_readra;         // nios2_0_custom_instruction_master_multi_xconnect:ci_master1_readra -> nios2_0_custom_instruction_master_multi_slave_translator1:ci_slave_readra
	wire   [4:0] nios2_0_custom_instruction_master_multi_xconnect_ci_master1_a;              // nios2_0_custom_instruction_master_multi_xconnect:ci_master1_a -> nios2_0_custom_instruction_master_multi_slave_translator1:ci_slave_a
	wire   [4:0] nios2_0_custom_instruction_master_multi_xconnect_ci_master1_b;              // nios2_0_custom_instruction_master_multi_xconnect:ci_master1_b -> nios2_0_custom_instruction_master_multi_slave_translator1:ci_slave_b
	wire         nios2_0_custom_instruction_master_multi_xconnect_ci_master1_readrb;         // nios2_0_custom_instruction_master_multi_xconnect:ci_master1_readrb -> nios2_0_custom_instruction_master_multi_slave_translator1:ci_slave_readrb
	wire   [4:0] nios2_0_custom_instruction_master_multi_xconnect_ci_master1_c;              // nios2_0_custom_instruction_master_multi_xconnect:ci_master1_c -> nios2_0_custom_instruction_master_multi_slave_translator1:ci_slave_c
	wire         nios2_0_custom_instruction_master_multi_xconnect_ci_master1_clk;            // nios2_0_custom_instruction_master_multi_xconnect:ci_master1_clk -> nios2_0_custom_instruction_master_multi_slave_translator1:ci_slave_clk
	wire  [31:0] nios2_0_custom_instruction_master_multi_xconnect_ci_master1_ipending;       // nios2_0_custom_instruction_master_multi_xconnect:ci_master1_ipending -> nios2_0_custom_instruction_master_multi_slave_translator1:ci_slave_ipending
	wire         nios2_0_custom_instruction_master_multi_xconnect_ci_master1_start;          // nios2_0_custom_instruction_master_multi_xconnect:ci_master1_start -> nios2_0_custom_instruction_master_multi_slave_translator1:ci_slave_start
	wire         nios2_0_custom_instruction_master_multi_xconnect_ci_master1_reset_req;      // nios2_0_custom_instruction_master_multi_xconnect:ci_master1_reset_req -> nios2_0_custom_instruction_master_multi_slave_translator1:ci_slave_reset_req
	wire         nios2_0_custom_instruction_master_multi_xconnect_ci_master1_done;           // nios2_0_custom_instruction_master_multi_slave_translator1:ci_slave_done -> nios2_0_custom_instruction_master_multi_xconnect:ci_master1_done
	wire   [7:0] nios2_0_custom_instruction_master_multi_xconnect_ci_master1_n;              // nios2_0_custom_instruction_master_multi_xconnect:ci_master1_n -> nios2_0_custom_instruction_master_multi_slave_translator1:ci_slave_n
	wire  [31:0] nios2_0_custom_instruction_master_multi_xconnect_ci_master1_result;         // nios2_0_custom_instruction_master_multi_slave_translator1:ci_slave_result -> nios2_0_custom_instruction_master_multi_xconnect:ci_master1_result
	wire         nios2_0_custom_instruction_master_multi_xconnect_ci_master1_estatus;        // nios2_0_custom_instruction_master_multi_xconnect:ci_master1_estatus -> nios2_0_custom_instruction_master_multi_slave_translator1:ci_slave_estatus
	wire         nios2_0_custom_instruction_master_multi_xconnect_ci_master1_clk_en;         // nios2_0_custom_instruction_master_multi_xconnect:ci_master1_clken -> nios2_0_custom_instruction_master_multi_slave_translator1:ci_slave_clken
	wire  [31:0] nios2_0_custom_instruction_master_multi_xconnect_ci_master1_datab;          // nios2_0_custom_instruction_master_multi_xconnect:ci_master1_datab -> nios2_0_custom_instruction_master_multi_slave_translator1:ci_slave_datab
	wire  [31:0] nios2_0_custom_instruction_master_multi_xconnect_ci_master1_dataa;          // nios2_0_custom_instruction_master_multi_xconnect:ci_master1_dataa -> nios2_0_custom_instruction_master_multi_slave_translator1:ci_slave_dataa
	wire         nios2_0_custom_instruction_master_multi_xconnect_ci_master1_reset;          // nios2_0_custom_instruction_master_multi_xconnect:ci_master1_reset -> nios2_0_custom_instruction_master_multi_slave_translator1:ci_slave_reset
	wire         nios2_0_custom_instruction_master_multi_xconnect_ci_master1_writerc;        // nios2_0_custom_instruction_master_multi_xconnect:ci_master1_writerc -> nios2_0_custom_instruction_master_multi_slave_translator1:ci_slave_writerc
	wire  [31:0] nios2_0_custom_instruction_master_multi_slave_translator1_ci_master_result; // acc_recv_0:result -> nios2_0_custom_instruction_master_multi_slave_translator1:ci_master_result
	wire         nios2_0_custom_instruction_master_multi_slave_translator1_ci_master_clk;    // nios2_0_custom_instruction_master_multi_slave_translator1:ci_master_clk -> acc_recv_0:nios_clk
	wire         nios2_0_custom_instruction_master_multi_slave_translator1_ci_master_clk_en; // nios2_0_custom_instruction_master_multi_slave_translator1:ci_master_clken -> acc_recv_0:clk_en
	wire  [31:0] nios2_0_custom_instruction_master_multi_slave_translator1_ci_master_datab;  // nios2_0_custom_instruction_master_multi_slave_translator1:ci_master_datab -> acc_recv_0:data_in_b
	wire  [31:0] nios2_0_custom_instruction_master_multi_slave_translator1_ci_master_dataa;  // nios2_0_custom_instruction_master_multi_slave_translator1:ci_master_dataa -> acc_recv_0:data_in_a
	wire         nios2_0_custom_instruction_master_multi_slave_translator1_ci_master_start;  // nios2_0_custom_instruction_master_multi_slave_translator1:ci_master_start -> acc_recv_0:start
	wire         nios2_0_custom_instruction_master_multi_slave_translator1_ci_master_reset;  // nios2_0_custom_instruction_master_multi_slave_translator1:ci_master_reset -> acc_recv_0:reset
	wire         nios2_0_custom_instruction_master_multi_slave_translator1_ci_master_done;   // acc_recv_0:done -> nios2_0_custom_instruction_master_multi_slave_translator1:ci_master_done
	wire   [2:0] nios2_0_custom_instruction_master_multi_slave_translator1_ci_master_n;      // nios2_0_custom_instruction_master_multi_slave_translator1:ci_master_n -> acc_recv_0:in_opcode
	wire         arbit_0_avalon_master_chipselect;                                           // arbit_0:chipselect -> mm_interconnect_0:arbit_0_avalon_master_chipselect
	wire         arbit_0_avalon_master_waitrequest;                                          // mm_interconnect_0:arbit_0_avalon_master_waitrequest -> arbit_0:waitrequest
	wire  [31:0] arbit_0_avalon_master_readdata;                                             // mm_interconnect_0:arbit_0_avalon_master_readdata -> arbit_0:readdata
	wire         arbit_0_avalon_master_read;                                                 // arbit_0:read -> mm_interconnect_0:arbit_0_avalon_master_read
	wire  [19:0] arbit_0_avalon_master_address;                                              // arbit_0:mem_addr -> mm_interconnect_0:arbit_0_avalon_master_address
	wire  [31:0] arbit_0_avalon_master_writedata;                                            // arbit_0:writedata -> mm_interconnect_0:arbit_0_avalon_master_writedata
	wire         arbit_0_avalon_master_write;                                                // arbit_0:write -> mm_interconnect_0:arbit_0_avalon_master_write
	wire         mm_interconnect_0_mem_s2_chipselect;                                        // mm_interconnect_0:mem_s2_chipselect -> mem:chipselect2
	wire  [31:0] mm_interconnect_0_mem_s2_readdata;                                          // mem:readdata2 -> mm_interconnect_0:mem_s2_readdata
	wire  [17:0] mm_interconnect_0_mem_s2_address;                                           // mm_interconnect_0:mem_s2_address -> mem:address2
	wire   [3:0] mm_interconnect_0_mem_s2_byteenable;                                        // mm_interconnect_0:mem_s2_byteenable -> mem:byteenable2
	wire         mm_interconnect_0_mem_s2_write;                                             // mm_interconnect_0:mem_s2_write -> mem:write2
	wire  [31:0] mm_interconnect_0_mem_s2_writedata;                                         // mm_interconnect_0:mem_s2_writedata -> mem:writedata2
	wire         mm_interconnect_0_mem_s2_clken;                                             // mm_interconnect_0:mem_s2_clken -> mem:clken2
	wire  [31:0] nios2_0_data_master_readdata;                                               // mm_interconnect_1:nios2_0_data_master_readdata -> nios2_0:d_readdata
	wire         nios2_0_data_master_waitrequest;                                            // mm_interconnect_1:nios2_0_data_master_waitrequest -> nios2_0:d_waitrequest
	wire         nios2_0_data_master_debugaccess;                                            // nios2_0:debug_mem_slave_debugaccess_to_roms -> mm_interconnect_1:nios2_0_data_master_debugaccess
	wire  [20:0] nios2_0_data_master_address;                                                // nios2_0:d_address -> mm_interconnect_1:nios2_0_data_master_address
	wire   [3:0] nios2_0_data_master_byteenable;                                             // nios2_0:d_byteenable -> mm_interconnect_1:nios2_0_data_master_byteenable
	wire         nios2_0_data_master_read;                                                   // nios2_0:d_read -> mm_interconnect_1:nios2_0_data_master_read
	wire         nios2_0_data_master_readdatavalid;                                          // mm_interconnect_1:nios2_0_data_master_readdatavalid -> nios2_0:d_readdatavalid
	wire         nios2_0_data_master_write;                                                  // nios2_0:d_write -> mm_interconnect_1:nios2_0_data_master_write
	wire  [31:0] nios2_0_data_master_writedata;                                              // nios2_0:d_writedata -> mm_interconnect_1:nios2_0_data_master_writedata
	wire  [31:0] nios2_0_instruction_master_readdata;                                        // mm_interconnect_1:nios2_0_instruction_master_readdata -> nios2_0:i_readdata
	wire         nios2_0_instruction_master_waitrequest;                                     // mm_interconnect_1:nios2_0_instruction_master_waitrequest -> nios2_0:i_waitrequest
	wire  [20:0] nios2_0_instruction_master_address;                                         // nios2_0:i_address -> mm_interconnect_1:nios2_0_instruction_master_address
	wire         nios2_0_instruction_master_read;                                            // nios2_0:i_read -> mm_interconnect_1:nios2_0_instruction_master_read
	wire         nios2_0_instruction_master_readdatavalid;                                   // mm_interconnect_1:nios2_0_instruction_master_readdatavalid -> nios2_0:i_readdatavalid
	wire         mm_interconnect_1_jtaguart_0_avalon_jtag_slave_chipselect;                  // mm_interconnect_1:jtaguart_0_avalon_jtag_slave_chipselect -> jtaguart_0:av_chipselect
	wire  [31:0] mm_interconnect_1_jtaguart_0_avalon_jtag_slave_readdata;                    // jtaguart_0:av_readdata -> mm_interconnect_1:jtaguart_0_avalon_jtag_slave_readdata
	wire         mm_interconnect_1_jtaguart_0_avalon_jtag_slave_waitrequest;                 // jtaguart_0:av_waitrequest -> mm_interconnect_1:jtaguart_0_avalon_jtag_slave_waitrequest
	wire   [0:0] mm_interconnect_1_jtaguart_0_avalon_jtag_slave_address;                     // mm_interconnect_1:jtaguart_0_avalon_jtag_slave_address -> jtaguart_0:av_address
	wire         mm_interconnect_1_jtaguart_0_avalon_jtag_slave_read;                        // mm_interconnect_1:jtaguart_0_avalon_jtag_slave_read -> jtaguart_0:av_read_n
	wire         mm_interconnect_1_jtaguart_0_avalon_jtag_slave_write;                       // mm_interconnect_1:jtaguart_0_avalon_jtag_slave_write -> jtaguart_0:av_write_n
	wire  [31:0] mm_interconnect_1_jtaguart_0_avalon_jtag_slave_writedata;                   // mm_interconnect_1:jtaguart_0_avalon_jtag_slave_writedata -> jtaguart_0:av_writedata
	wire  [31:0] mm_interconnect_1_sysid_control_slave_readdata;                             // sysid:readdata -> mm_interconnect_1:sysid_control_slave_readdata
	wire   [0:0] mm_interconnect_1_sysid_control_slave_address;                              // mm_interconnect_1:sysid_control_slave_address -> sysid:address
	wire  [31:0] mm_interconnect_1_performance_counter_0_control_slave_readdata;             // performance_counter_0:readdata -> mm_interconnect_1:performance_counter_0_control_slave_readdata
	wire   [3:0] mm_interconnect_1_performance_counter_0_control_slave_address;              // mm_interconnect_1:performance_counter_0_control_slave_address -> performance_counter_0:address
	wire         mm_interconnect_1_performance_counter_0_control_slave_begintransfer;        // mm_interconnect_1:performance_counter_0_control_slave_begintransfer -> performance_counter_0:begintransfer
	wire         mm_interconnect_1_performance_counter_0_control_slave_write;                // mm_interconnect_1:performance_counter_0_control_slave_write -> performance_counter_0:write
	wire  [31:0] mm_interconnect_1_performance_counter_0_control_slave_writedata;            // mm_interconnect_1:performance_counter_0_control_slave_writedata -> performance_counter_0:writedata
	wire  [31:0] mm_interconnect_1_nios2_0_debug_mem_slave_readdata;                         // nios2_0:debug_mem_slave_readdata -> mm_interconnect_1:nios2_0_debug_mem_slave_readdata
	wire         mm_interconnect_1_nios2_0_debug_mem_slave_waitrequest;                      // nios2_0:debug_mem_slave_waitrequest -> mm_interconnect_1:nios2_0_debug_mem_slave_waitrequest
	wire         mm_interconnect_1_nios2_0_debug_mem_slave_debugaccess;                      // mm_interconnect_1:nios2_0_debug_mem_slave_debugaccess -> nios2_0:debug_mem_slave_debugaccess
	wire   [8:0] mm_interconnect_1_nios2_0_debug_mem_slave_address;                          // mm_interconnect_1:nios2_0_debug_mem_slave_address -> nios2_0:debug_mem_slave_address
	wire         mm_interconnect_1_nios2_0_debug_mem_slave_read;                             // mm_interconnect_1:nios2_0_debug_mem_slave_read -> nios2_0:debug_mem_slave_read
	wire   [3:0] mm_interconnect_1_nios2_0_debug_mem_slave_byteenable;                       // mm_interconnect_1:nios2_0_debug_mem_slave_byteenable -> nios2_0:debug_mem_slave_byteenable
	wire         mm_interconnect_1_nios2_0_debug_mem_slave_write;                            // mm_interconnect_1:nios2_0_debug_mem_slave_write -> nios2_0:debug_mem_slave_write
	wire  [31:0] mm_interconnect_1_nios2_0_debug_mem_slave_writedata;                        // mm_interconnect_1:nios2_0_debug_mem_slave_writedata -> nios2_0:debug_mem_slave_writedata
	wire         mm_interconnect_1_sys_clk_timer_s1_chipselect;                              // mm_interconnect_1:sys_clk_timer_s1_chipselect -> sys_clk_timer:chipselect
	wire  [15:0] mm_interconnect_1_sys_clk_timer_s1_readdata;                                // sys_clk_timer:readdata -> mm_interconnect_1:sys_clk_timer_s1_readdata
	wire   [2:0] mm_interconnect_1_sys_clk_timer_s1_address;                                 // mm_interconnect_1:sys_clk_timer_s1_address -> sys_clk_timer:address
	wire         mm_interconnect_1_sys_clk_timer_s1_write;                                   // mm_interconnect_1:sys_clk_timer_s1_write -> sys_clk_timer:write_n
	wire  [15:0] mm_interconnect_1_sys_clk_timer_s1_writedata;                               // mm_interconnect_1:sys_clk_timer_s1_writedata -> sys_clk_timer:writedata
	wire         mm_interconnect_1_mem_s1_chipselect;                                        // mm_interconnect_1:mem_s1_chipselect -> mem:chipselect
	wire  [31:0] mm_interconnect_1_mem_s1_readdata;                                          // mem:readdata -> mm_interconnect_1:mem_s1_readdata
	wire  [17:0] mm_interconnect_1_mem_s1_address;                                           // mm_interconnect_1:mem_s1_address -> mem:address
	wire   [3:0] mm_interconnect_1_mem_s1_byteenable;                                        // mm_interconnect_1:mem_s1_byteenable -> mem:byteenable
	wire         mm_interconnect_1_mem_s1_write;                                             // mm_interconnect_1:mem_s1_write -> mem:write
	wire  [31:0] mm_interconnect_1_mem_s1_writedata;                                         // mm_interconnect_1:mem_s1_writedata -> mem:writedata
	wire         mm_interconnect_1_mem_s1_clken;                                             // mm_interconnect_1:mem_s1_clken -> mem:clken
	wire         irq_mapper_receiver0_irq;                                                   // sys_clk_timer:irq -> irq_mapper:receiver0_irq
	wire         irq_mapper_receiver1_irq;                                                   // jtaguart_0:av_irq -> irq_mapper:receiver1_irq
	wire  [31:0] nios2_0_irq_irq;                                                            // irq_mapper:sender_irq -> nios2_0:irq
	wire         rst_controller_reset_out_reset;                                             // rst_controller:reset_out -> [arbit_0:reset, irq_mapper:reset, jtaguart_0:rst_n, mem:reset, mem:reset2, mm_interconnect_0:arbit_0_reset_reset_bridge_in_reset_reset, mm_interconnect_1:nios2_0_reset_reset_bridge_in_reset_reset, nios2_0:reset_n, performance_counter_0:reset_n, rst_translator:in_reset, sys_clk_timer:reset_n, sysid:reset_n]
	wire         rst_controller_reset_out_reset_req;                                         // rst_controller:reset_req -> [mem:reset_req, mem:reset_req2, nios2_0:reset_req, rst_translator:reset_req_in]

	acc_send #(
		.cpu_width        (32),
		.packetizer_width (128),
		.data_width       (32),
		.mem_width        (32),
		.mem_depth        (11),
		.threshold        (1),
		.SIZE             (3)
	) acc_0 (
		.packet           (acc_0_packet_out_packet),                                                    //                      packet_out.packet
		.packet_out_valid (acc_0_packet_out_valid),                                                     //                                .valid
		.data_in_a        (nios2_0_custom_instruction_master_multi_slave_translator0_ci_master_dataa),  // nios_custom_instruction_slave_1.dataa
		.data_in_b        (nios2_0_custom_instruction_master_multi_slave_translator0_ci_master_datab),  //                                .datab
		.in_opcode        (nios2_0_custom_instruction_master_multi_slave_translator0_ci_master_n),      //                                .n
		.start            (nios2_0_custom_instruction_master_multi_slave_translator0_ci_master_start),  //                                .start
		.result           (nios2_0_custom_instruction_master_multi_slave_translator0_ci_master_result), //                                .result
		.done             (nios2_0_custom_instruction_master_multi_slave_translator0_ci_master_done),   //                                .done
		.nios_clk         (nios2_0_custom_instruction_master_multi_slave_translator0_ci_master_clk),    //                                .clk
		.reset            (nios2_0_custom_instruction_master_multi_slave_translator0_ci_master_reset),  //                                .reset
		.clk_en           (nios2_0_custom_instruction_master_multi_slave_translator0_ci_master_clk_en)  //                                .clk_en
	);

	acc_recv #(
		.cpu_width        (32),
		.packetizer_width (128),
		.data_width       (32),
		.CONTENT_WIDTH    (36),
		.mem_width        (32),
		.mem_depth        (11),
		.threshold        (1),
		.SIZE             (3)
	) acc_recv_0 (
		.packet_in       (acc_recv_0_pack_in_packet),                                                  //                         pack_in.packet
		.packet_in_valid (acc_recv_0_pack_in_valid),                                                   //                                .valid
		.nios_clk        (nios2_0_custom_instruction_master_multi_slave_translator1_ci_master_clk),    // nios_custom_instruction_slave_2.clk
		.clk_en          (nios2_0_custom_instruction_master_multi_slave_translator1_ci_master_clk_en), //                                .clk_en
		.data_in_a       (nios2_0_custom_instruction_master_multi_slave_translator1_ci_master_dataa),  //                                .dataa
		.data_in_b       (nios2_0_custom_instruction_master_multi_slave_translator1_ci_master_datab),  //                                .datab
		.in_opcode       (nios2_0_custom_instruction_master_multi_slave_translator1_ci_master_n),      //                                .n
		.start           (nios2_0_custom_instruction_master_multi_slave_translator1_ci_master_start),  //                                .start
		.result          (nios2_0_custom_instruction_master_multi_slave_translator1_ci_master_result), //                                .result
		.done            (nios2_0_custom_instruction_master_multi_slave_translator1_ci_master_done),   //                                .done
		.reset           (nios2_0_custom_instruction_master_multi_slave_translator1_ci_master_reset),  //                                .reset
		.data_to_mem     (acc_recv_0_conduit_end_data_to_mem),                                         //                     conduit_end.data_to_mem
		.write           (acc_recv_0_conduit_end_write),                                               //                                .write
		.write_addr      (acc_recv_0_conduit_end_write_addr)                                           //                                .write_addr
	);

	arbit #(
		.cpu_width        (32),
		.packetizer_width (128),
		.data_width       (32),
		.mem_width        (32),
		.mem_depth        (11),
		.threshold        (1),
		.SIZE             (3)
	) arbit_0 (
		.chipselect    (arbit_0_avalon_master_chipselect),   // avalon_master.chipselect
		.writedata     (arbit_0_avalon_master_writedata),    //              .writedata
		.waitrequest   (arbit_0_avalon_master_waitrequest),  //              .waitrequest
		.write         (arbit_0_avalon_master_write),        //              .write
		.read          (arbit_0_avalon_master_read),         //              .read
		.readdata      (arbit_0_avalon_master_readdata),     //              .readdata
		.mem_addr      (arbit_0_avalon_master_address),      //              .address
		.write_addr_r  (acc_recv_0_conduit_end_write_addr),  //         acc_r.write_addr
		.write_r       (acc_recv_0_conduit_end_write),       //              .write
		.data_to_mem_r (acc_recv_0_conduit_end_data_to_mem), //              .data_to_mem
		.clk           (pll_0_outclk0_clk),                  //         clock.clk
		.reset         (rst_controller_reset_out_reset)      //         reset.reset
	);

	nios2_jtaguart_0 jtaguart_0 (
		.clk            (pll_0_outclk0_clk),                                          //               clk.clk
		.rst_n          (~rst_controller_reset_out_reset),                            //             reset.reset_n
		.av_chipselect  (mm_interconnect_1_jtaguart_0_avalon_jtag_slave_chipselect),  // avalon_jtag_slave.chipselect
		.av_address     (mm_interconnect_1_jtaguart_0_avalon_jtag_slave_address),     //                  .address
		.av_read_n      (~mm_interconnect_1_jtaguart_0_avalon_jtag_slave_read),       //                  .read_n
		.av_readdata    (mm_interconnect_1_jtaguart_0_avalon_jtag_slave_readdata),    //                  .readdata
		.av_write_n     (~mm_interconnect_1_jtaguart_0_avalon_jtag_slave_write),      //                  .write_n
		.av_writedata   (mm_interconnect_1_jtaguart_0_avalon_jtag_slave_writedata),   //                  .writedata
		.av_waitrequest (mm_interconnect_1_jtaguart_0_avalon_jtag_slave_waitrequest), //                  .waitrequest
		.av_irq         (irq_mapper_receiver1_irq)                                    //               irq.irq
	);

	nios2_mem mem (
		.clk         (pll_0_outclk0_clk),                   //   clk1.clk
		.address     (mm_interconnect_1_mem_s1_address),    //     s1.address
		.clken       (mm_interconnect_1_mem_s1_clken),      //       .clken
		.chipselect  (mm_interconnect_1_mem_s1_chipselect), //       .chipselect
		.write       (mm_interconnect_1_mem_s1_write),      //       .write
		.readdata    (mm_interconnect_1_mem_s1_readdata),   //       .readdata
		.writedata   (mm_interconnect_1_mem_s1_writedata),  //       .writedata
		.byteenable  (mm_interconnect_1_mem_s1_byteenable), //       .byteenable
		.reset       (rst_controller_reset_out_reset),      // reset1.reset
		.reset_req   (rst_controller_reset_out_reset_req),  //       .reset_req
		.address2    (mm_interconnect_0_mem_s2_address),    //     s2.address
		.chipselect2 (mm_interconnect_0_mem_s2_chipselect), //       .chipselect
		.clken2      (mm_interconnect_0_mem_s2_clken),      //       .clken
		.write2      (mm_interconnect_0_mem_s2_write),      //       .write
		.readdata2   (mm_interconnect_0_mem_s2_readdata),   //       .readdata
		.writedata2  (mm_interconnect_0_mem_s2_writedata),  //       .writedata
		.byteenable2 (mm_interconnect_0_mem_s2_byteenable), //       .byteenable
		.clk2        (pll_0_outclk0_clk),                   //   clk2.clk
		.reset2      (rst_controller_reset_out_reset),      // reset2.reset
		.reset_req2  (rst_controller_reset_out_reset_req)   //       .reset_req
	);

	nios2_nios2_0 nios2_0 (
		.clk                                 (pll_0_outclk0_clk),                                     //                       clk.clk
		.reset_n                             (~rst_controller_reset_out_reset),                       //                     reset.reset_n
		.reset_req                           (rst_controller_reset_out_reset_req),                    //                          .reset_req
		.d_address                           (nios2_0_data_master_address),                           //               data_master.address
		.d_byteenable                        (nios2_0_data_master_byteenable),                        //                          .byteenable
		.d_read                              (nios2_0_data_master_read),                              //                          .read
		.d_readdata                          (nios2_0_data_master_readdata),                          //                          .readdata
		.d_waitrequest                       (nios2_0_data_master_waitrequest),                       //                          .waitrequest
		.d_write                             (nios2_0_data_master_write),                             //                          .write
		.d_writedata                         (nios2_0_data_master_writedata),                         //                          .writedata
		.d_readdatavalid                     (nios2_0_data_master_readdatavalid),                     //                          .readdatavalid
		.debug_mem_slave_debugaccess_to_roms (nios2_0_data_master_debugaccess),                       //                          .debugaccess
		.i_address                           (nios2_0_instruction_master_address),                    //        instruction_master.address
		.i_read                              (nios2_0_instruction_master_read),                       //                          .read
		.i_readdata                          (nios2_0_instruction_master_readdata),                   //                          .readdata
		.i_waitrequest                       (nios2_0_instruction_master_waitrequest),                //                          .waitrequest
		.i_readdatavalid                     (nios2_0_instruction_master_readdatavalid),              //                          .readdatavalid
		.irq                                 (nios2_0_irq_irq),                                       //                       irq.irq
		.debug_reset_request                 (),                                                      //       debug_reset_request.reset
		.debug_mem_slave_address             (mm_interconnect_1_nios2_0_debug_mem_slave_address),     //           debug_mem_slave.address
		.debug_mem_slave_byteenable          (mm_interconnect_1_nios2_0_debug_mem_slave_byteenable),  //                          .byteenable
		.debug_mem_slave_debugaccess         (mm_interconnect_1_nios2_0_debug_mem_slave_debugaccess), //                          .debugaccess
		.debug_mem_slave_read                (mm_interconnect_1_nios2_0_debug_mem_slave_read),        //                          .read
		.debug_mem_slave_readdata            (mm_interconnect_1_nios2_0_debug_mem_slave_readdata),    //                          .readdata
		.debug_mem_slave_waitrequest         (mm_interconnect_1_nios2_0_debug_mem_slave_waitrequest), //                          .waitrequest
		.debug_mem_slave_write               (mm_interconnect_1_nios2_0_debug_mem_slave_write),       //                          .write
		.debug_mem_slave_writedata           (mm_interconnect_1_nios2_0_debug_mem_slave_writedata),   //                          .writedata
		.A_ci_multi_done                     (nios2_0_custom_instruction_master_done),                // custom_instruction_master.done
		.A_ci_multi_result                   (nios2_0_custom_instruction_master_multi_result),        //                          .multi_result
		.A_ci_multi_a                        (nios2_0_custom_instruction_master_multi_a),             //                          .multi_a
		.A_ci_multi_b                        (nios2_0_custom_instruction_master_multi_b),             //                          .multi_b
		.A_ci_multi_c                        (nios2_0_custom_instruction_master_multi_c),             //                          .multi_c
		.A_ci_multi_clk_en                   (nios2_0_custom_instruction_master_clk_en),              //                          .clk_en
		.A_ci_multi_clock                    (nios2_0_custom_instruction_master_clk),                 //                          .clk
		.A_ci_multi_reset                    (nios2_0_custom_instruction_master_reset),               //                          .reset
		.A_ci_multi_reset_req                (nios2_0_custom_instruction_master_reset_req),           //                          .reset_req
		.A_ci_multi_dataa                    (nios2_0_custom_instruction_master_multi_dataa),         //                          .multi_dataa
		.A_ci_multi_datab                    (nios2_0_custom_instruction_master_multi_datab),         //                          .multi_datab
		.A_ci_multi_n                        (nios2_0_custom_instruction_master_multi_n),             //                          .multi_n
		.A_ci_multi_readra                   (nios2_0_custom_instruction_master_multi_readra),        //                          .multi_readra
		.A_ci_multi_readrb                   (nios2_0_custom_instruction_master_multi_readrb),        //                          .multi_readrb
		.A_ci_multi_start                    (nios2_0_custom_instruction_master_start),               //                          .start
		.A_ci_multi_writerc                  (nios2_0_custom_instruction_master_multi_writerc)        //                          .multi_writerc
	);

	nios2_performance_counter_0 performance_counter_0 (
		.clk           (pll_0_outclk0_clk),                                                   //           clk.clk
		.reset_n       (~rst_controller_reset_out_reset),                                     //         reset.reset_n
		.address       (mm_interconnect_1_performance_counter_0_control_slave_address),       // control_slave.address
		.begintransfer (mm_interconnect_1_performance_counter_0_control_slave_begintransfer), //              .begintransfer
		.readdata      (mm_interconnect_1_performance_counter_0_control_slave_readdata),      //              .readdata
		.write         (mm_interconnect_1_performance_counter_0_control_slave_write),         //              .write
		.writedata     (mm_interconnect_1_performance_counter_0_control_slave_writedata)      //              .writedata
	);

	nios2_pll_0 pll_0 (
		.refclk   (clk_clk),           //  refclk.clk
		.rst      (~reset_reset_n),    //   reset.reset
		.outclk_0 (pll_0_outclk0_clk), // outclk0.clk
		.locked   ()                   // (terminated)
	);

	nios2_sys_clk_timer sys_clk_timer (
		.clk        (pll_0_outclk0_clk),                             //   clk.clk
		.reset_n    (~rst_controller_reset_out_reset),               // reset.reset_n
		.address    (mm_interconnect_1_sys_clk_timer_s1_address),    //    s1.address
		.writedata  (mm_interconnect_1_sys_clk_timer_s1_writedata),  //      .writedata
		.readdata   (mm_interconnect_1_sys_clk_timer_s1_readdata),   //      .readdata
		.chipselect (mm_interconnect_1_sys_clk_timer_s1_chipselect), //      .chipselect
		.write_n    (~mm_interconnect_1_sys_clk_timer_s1_write),     //      .write_n
		.irq        (irq_mapper_receiver0_irq)                       //   irq.irq
	);

	nios2_sysid sysid (
		.clock    (pll_0_outclk0_clk),                              //           clk.clk
		.reset_n  (~rst_controller_reset_out_reset),                //         reset.reset_n
		.readdata (mm_interconnect_1_sysid_control_slave_readdata), // control_slave.readdata
		.address  (mm_interconnect_1_sysid_control_slave_address)   //              .address
	);

	altera_customins_master_translator #(
		.SHARED_COMB_AND_MULTI (0)
	) nios2_0_custom_instruction_master_translator (
		.ci_slave_result           (),                                                                       //        ci_slave.result
		.ci_slave_multi_clk        (nios2_0_custom_instruction_master_clk),                                  //                .clk
		.ci_slave_multi_reset      (nios2_0_custom_instruction_master_reset),                                //                .reset
		.ci_slave_multi_clken      (nios2_0_custom_instruction_master_clk_en),                               //                .clk_en
		.ci_slave_multi_reset_req  (nios2_0_custom_instruction_master_reset_req),                            //                .reset_req
		.ci_slave_multi_start      (nios2_0_custom_instruction_master_start),                                //                .start
		.ci_slave_multi_done       (nios2_0_custom_instruction_master_done),                                 //                .done
		.ci_slave_multi_dataa      (nios2_0_custom_instruction_master_multi_dataa),                          //                .multi_dataa
		.ci_slave_multi_datab      (nios2_0_custom_instruction_master_multi_datab),                          //                .multi_datab
		.ci_slave_multi_result     (nios2_0_custom_instruction_master_multi_result),                         //                .multi_result
		.ci_slave_multi_n          (nios2_0_custom_instruction_master_multi_n),                              //                .multi_n
		.ci_slave_multi_readra     (nios2_0_custom_instruction_master_multi_readra),                         //                .multi_readra
		.ci_slave_multi_readrb     (nios2_0_custom_instruction_master_multi_readrb),                         //                .multi_readrb
		.ci_slave_multi_writerc    (nios2_0_custom_instruction_master_multi_writerc),                        //                .multi_writerc
		.ci_slave_multi_a          (nios2_0_custom_instruction_master_multi_a),                              //                .multi_a
		.ci_slave_multi_b          (nios2_0_custom_instruction_master_multi_b),                              //                .multi_b
		.ci_slave_multi_c          (nios2_0_custom_instruction_master_multi_c),                              //                .multi_c
		.comb_ci_master_result     (),                                                                       //  comb_ci_master.result
		.multi_ci_master_clk       (nios2_0_custom_instruction_master_translator_multi_ci_master_clk),       // multi_ci_master.clk
		.multi_ci_master_reset     (nios2_0_custom_instruction_master_translator_multi_ci_master_reset),     //                .reset
		.multi_ci_master_clken     (nios2_0_custom_instruction_master_translator_multi_ci_master_clk_en),    //                .clk_en
		.multi_ci_master_reset_req (nios2_0_custom_instruction_master_translator_multi_ci_master_reset_req), //                .reset_req
		.multi_ci_master_start     (nios2_0_custom_instruction_master_translator_multi_ci_master_start),     //                .start
		.multi_ci_master_done      (nios2_0_custom_instruction_master_translator_multi_ci_master_done),      //                .done
		.multi_ci_master_dataa     (nios2_0_custom_instruction_master_translator_multi_ci_master_dataa),     //                .dataa
		.multi_ci_master_datab     (nios2_0_custom_instruction_master_translator_multi_ci_master_datab),     //                .datab
		.multi_ci_master_result    (nios2_0_custom_instruction_master_translator_multi_ci_master_result),    //                .result
		.multi_ci_master_n         (nios2_0_custom_instruction_master_translator_multi_ci_master_n),         //                .n
		.multi_ci_master_readra    (nios2_0_custom_instruction_master_translator_multi_ci_master_readra),    //                .readra
		.multi_ci_master_readrb    (nios2_0_custom_instruction_master_translator_multi_ci_master_readrb),    //                .readrb
		.multi_ci_master_writerc   (nios2_0_custom_instruction_master_translator_multi_ci_master_writerc),   //                .writerc
		.multi_ci_master_a         (nios2_0_custom_instruction_master_translator_multi_ci_master_a),         //                .a
		.multi_ci_master_b         (nios2_0_custom_instruction_master_translator_multi_ci_master_b),         //                .b
		.multi_ci_master_c         (nios2_0_custom_instruction_master_translator_multi_ci_master_c),         //                .c
		.ci_slave_dataa            (32'b00000000000000000000000000000000),                                   //     (terminated)
		.ci_slave_datab            (32'b00000000000000000000000000000000),                                   //     (terminated)
		.ci_slave_n                (8'b00000000),                                                            //     (terminated)
		.ci_slave_readra           (1'b0),                                                                   //     (terminated)
		.ci_slave_readrb           (1'b0),                                                                   //     (terminated)
		.ci_slave_writerc          (1'b0),                                                                   //     (terminated)
		.ci_slave_a                (5'b00000),                                                               //     (terminated)
		.ci_slave_b                (5'b00000),                                                               //     (terminated)
		.ci_slave_c                (5'b00000),                                                               //     (terminated)
		.ci_slave_ipending         (32'b00000000000000000000000000000000),                                   //     (terminated)
		.ci_slave_estatus          (1'b0),                                                                   //     (terminated)
		.comb_ci_master_dataa      (),                                                                       //     (terminated)
		.comb_ci_master_datab      (),                                                                       //     (terminated)
		.comb_ci_master_n          (),                                                                       //     (terminated)
		.comb_ci_master_readra     (),                                                                       //     (terminated)
		.comb_ci_master_readrb     (),                                                                       //     (terminated)
		.comb_ci_master_writerc    (),                                                                       //     (terminated)
		.comb_ci_master_a          (),                                                                       //     (terminated)
		.comb_ci_master_b          (),                                                                       //     (terminated)
		.comb_ci_master_c          (),                                                                       //     (terminated)
		.comb_ci_master_ipending   (),                                                                       //     (terminated)
		.comb_ci_master_estatus    ()                                                                        //     (terminated)
	);

	nios2_nios2_0_custom_instruction_master_multi_xconnect nios2_0_custom_instruction_master_multi_xconnect (
		.ci_slave_dataa       (nios2_0_custom_instruction_master_translator_multi_ci_master_dataa),     //   ci_slave.dataa
		.ci_slave_datab       (nios2_0_custom_instruction_master_translator_multi_ci_master_datab),     //           .datab
		.ci_slave_result      (nios2_0_custom_instruction_master_translator_multi_ci_master_result),    //           .result
		.ci_slave_n           (nios2_0_custom_instruction_master_translator_multi_ci_master_n),         //           .n
		.ci_slave_readra      (nios2_0_custom_instruction_master_translator_multi_ci_master_readra),    //           .readra
		.ci_slave_readrb      (nios2_0_custom_instruction_master_translator_multi_ci_master_readrb),    //           .readrb
		.ci_slave_writerc     (nios2_0_custom_instruction_master_translator_multi_ci_master_writerc),   //           .writerc
		.ci_slave_a           (nios2_0_custom_instruction_master_translator_multi_ci_master_a),         //           .a
		.ci_slave_b           (nios2_0_custom_instruction_master_translator_multi_ci_master_b),         //           .b
		.ci_slave_c           (nios2_0_custom_instruction_master_translator_multi_ci_master_c),         //           .c
		.ci_slave_ipending    (),                                                                       //           .ipending
		.ci_slave_estatus     (),                                                                       //           .estatus
		.ci_slave_clk         (nios2_0_custom_instruction_master_translator_multi_ci_master_clk),       //           .clk
		.ci_slave_reset       (nios2_0_custom_instruction_master_translator_multi_ci_master_reset),     //           .reset
		.ci_slave_clken       (nios2_0_custom_instruction_master_translator_multi_ci_master_clk_en),    //           .clk_en
		.ci_slave_reset_req   (nios2_0_custom_instruction_master_translator_multi_ci_master_reset_req), //           .reset_req
		.ci_slave_start       (nios2_0_custom_instruction_master_translator_multi_ci_master_start),     //           .start
		.ci_slave_done        (nios2_0_custom_instruction_master_translator_multi_ci_master_done),      //           .done
		.ci_master0_dataa     (nios2_0_custom_instruction_master_multi_xconnect_ci_master0_dataa),      // ci_master0.dataa
		.ci_master0_datab     (nios2_0_custom_instruction_master_multi_xconnect_ci_master0_datab),      //           .datab
		.ci_master0_result    (nios2_0_custom_instruction_master_multi_xconnect_ci_master0_result),     //           .result
		.ci_master0_n         (nios2_0_custom_instruction_master_multi_xconnect_ci_master0_n),          //           .n
		.ci_master0_readra    (nios2_0_custom_instruction_master_multi_xconnect_ci_master0_readra),     //           .readra
		.ci_master0_readrb    (nios2_0_custom_instruction_master_multi_xconnect_ci_master0_readrb),     //           .readrb
		.ci_master0_writerc   (nios2_0_custom_instruction_master_multi_xconnect_ci_master0_writerc),    //           .writerc
		.ci_master0_a         (nios2_0_custom_instruction_master_multi_xconnect_ci_master0_a),          //           .a
		.ci_master0_b         (nios2_0_custom_instruction_master_multi_xconnect_ci_master0_b),          //           .b
		.ci_master0_c         (nios2_0_custom_instruction_master_multi_xconnect_ci_master0_c),          //           .c
		.ci_master0_ipending  (nios2_0_custom_instruction_master_multi_xconnect_ci_master0_ipending),   //           .ipending
		.ci_master0_estatus   (nios2_0_custom_instruction_master_multi_xconnect_ci_master0_estatus),    //           .estatus
		.ci_master0_clk       (nios2_0_custom_instruction_master_multi_xconnect_ci_master0_clk),        //           .clk
		.ci_master0_reset     (nios2_0_custom_instruction_master_multi_xconnect_ci_master0_reset),      //           .reset
		.ci_master0_clken     (nios2_0_custom_instruction_master_multi_xconnect_ci_master0_clk_en),     //           .clk_en
		.ci_master0_reset_req (nios2_0_custom_instruction_master_multi_xconnect_ci_master0_reset_req),  //           .reset_req
		.ci_master0_start     (nios2_0_custom_instruction_master_multi_xconnect_ci_master0_start),      //           .start
		.ci_master0_done      (nios2_0_custom_instruction_master_multi_xconnect_ci_master0_done),       //           .done
		.ci_master1_dataa     (nios2_0_custom_instruction_master_multi_xconnect_ci_master1_dataa),      // ci_master1.dataa
		.ci_master1_datab     (nios2_0_custom_instruction_master_multi_xconnect_ci_master1_datab),      //           .datab
		.ci_master1_result    (nios2_0_custom_instruction_master_multi_xconnect_ci_master1_result),     //           .result
		.ci_master1_n         (nios2_0_custom_instruction_master_multi_xconnect_ci_master1_n),          //           .n
		.ci_master1_readra    (nios2_0_custom_instruction_master_multi_xconnect_ci_master1_readra),     //           .readra
		.ci_master1_readrb    (nios2_0_custom_instruction_master_multi_xconnect_ci_master1_readrb),     //           .readrb
		.ci_master1_writerc   (nios2_0_custom_instruction_master_multi_xconnect_ci_master1_writerc),    //           .writerc
		.ci_master1_a         (nios2_0_custom_instruction_master_multi_xconnect_ci_master1_a),          //           .a
		.ci_master1_b         (nios2_0_custom_instruction_master_multi_xconnect_ci_master1_b),          //           .b
		.ci_master1_c         (nios2_0_custom_instruction_master_multi_xconnect_ci_master1_c),          //           .c
		.ci_master1_ipending  (nios2_0_custom_instruction_master_multi_xconnect_ci_master1_ipending),   //           .ipending
		.ci_master1_estatus   (nios2_0_custom_instruction_master_multi_xconnect_ci_master1_estatus),    //           .estatus
		.ci_master1_clk       (nios2_0_custom_instruction_master_multi_xconnect_ci_master1_clk),        //           .clk
		.ci_master1_reset     (nios2_0_custom_instruction_master_multi_xconnect_ci_master1_reset),      //           .reset
		.ci_master1_clken     (nios2_0_custom_instruction_master_multi_xconnect_ci_master1_clk_en),     //           .clk_en
		.ci_master1_reset_req (nios2_0_custom_instruction_master_multi_xconnect_ci_master1_reset_req),  //           .reset_req
		.ci_master1_start     (nios2_0_custom_instruction_master_multi_xconnect_ci_master1_start),      //           .start
		.ci_master1_done      (nios2_0_custom_instruction_master_multi_xconnect_ci_master1_done)        //           .done
	);

	altera_customins_slave_translator #(
		.N_WIDTH          (3),
		.USE_DONE         (1),
		.NUM_FIXED_CYCLES (0)
	) nios2_0_custom_instruction_master_multi_slave_translator0 (
		.ci_slave_dataa      (nios2_0_custom_instruction_master_multi_xconnect_ci_master0_dataa),          //  ci_slave.dataa
		.ci_slave_datab      (nios2_0_custom_instruction_master_multi_xconnect_ci_master0_datab),          //          .datab
		.ci_slave_result     (nios2_0_custom_instruction_master_multi_xconnect_ci_master0_result),         //          .result
		.ci_slave_n          (nios2_0_custom_instruction_master_multi_xconnect_ci_master0_n),              //          .n
		.ci_slave_readra     (nios2_0_custom_instruction_master_multi_xconnect_ci_master0_readra),         //          .readra
		.ci_slave_readrb     (nios2_0_custom_instruction_master_multi_xconnect_ci_master0_readrb),         //          .readrb
		.ci_slave_writerc    (nios2_0_custom_instruction_master_multi_xconnect_ci_master0_writerc),        //          .writerc
		.ci_slave_a          (nios2_0_custom_instruction_master_multi_xconnect_ci_master0_a),              //          .a
		.ci_slave_b          (nios2_0_custom_instruction_master_multi_xconnect_ci_master0_b),              //          .b
		.ci_slave_c          (nios2_0_custom_instruction_master_multi_xconnect_ci_master0_c),              //          .c
		.ci_slave_ipending   (nios2_0_custom_instruction_master_multi_xconnect_ci_master0_ipending),       //          .ipending
		.ci_slave_estatus    (nios2_0_custom_instruction_master_multi_xconnect_ci_master0_estatus),        //          .estatus
		.ci_slave_clk        (nios2_0_custom_instruction_master_multi_xconnect_ci_master0_clk),            //          .clk
		.ci_slave_clken      (nios2_0_custom_instruction_master_multi_xconnect_ci_master0_clk_en),         //          .clk_en
		.ci_slave_reset_req  (nios2_0_custom_instruction_master_multi_xconnect_ci_master0_reset_req),      //          .reset_req
		.ci_slave_reset      (nios2_0_custom_instruction_master_multi_xconnect_ci_master0_reset),          //          .reset
		.ci_slave_start      (nios2_0_custom_instruction_master_multi_xconnect_ci_master0_start),          //          .start
		.ci_slave_done       (nios2_0_custom_instruction_master_multi_xconnect_ci_master0_done),           //          .done
		.ci_master_dataa     (nios2_0_custom_instruction_master_multi_slave_translator0_ci_master_dataa),  // ci_master.dataa
		.ci_master_datab     (nios2_0_custom_instruction_master_multi_slave_translator0_ci_master_datab),  //          .datab
		.ci_master_result    (nios2_0_custom_instruction_master_multi_slave_translator0_ci_master_result), //          .result
		.ci_master_n         (nios2_0_custom_instruction_master_multi_slave_translator0_ci_master_n),      //          .n
		.ci_master_clk       (nios2_0_custom_instruction_master_multi_slave_translator0_ci_master_clk),    //          .clk
		.ci_master_clken     (nios2_0_custom_instruction_master_multi_slave_translator0_ci_master_clk_en), //          .clk_en
		.ci_master_reset     (nios2_0_custom_instruction_master_multi_slave_translator0_ci_master_reset),  //          .reset
		.ci_master_start     (nios2_0_custom_instruction_master_multi_slave_translator0_ci_master_start),  //          .start
		.ci_master_done      (nios2_0_custom_instruction_master_multi_slave_translator0_ci_master_done),   //          .done
		.ci_master_readra    (),                                                                           // (terminated)
		.ci_master_readrb    (),                                                                           // (terminated)
		.ci_master_writerc   (),                                                                           // (terminated)
		.ci_master_a         (),                                                                           // (terminated)
		.ci_master_b         (),                                                                           // (terminated)
		.ci_master_c         (),                                                                           // (terminated)
		.ci_master_ipending  (),                                                                           // (terminated)
		.ci_master_estatus   (),                                                                           // (terminated)
		.ci_master_reset_req ()                                                                            // (terminated)
	);

	altera_customins_slave_translator #(
		.N_WIDTH          (3),
		.USE_DONE         (1),
		.NUM_FIXED_CYCLES (0)
	) nios2_0_custom_instruction_master_multi_slave_translator1 (
		.ci_slave_dataa      (nios2_0_custom_instruction_master_multi_xconnect_ci_master1_dataa),          //  ci_slave.dataa
		.ci_slave_datab      (nios2_0_custom_instruction_master_multi_xconnect_ci_master1_datab),          //          .datab
		.ci_slave_result     (nios2_0_custom_instruction_master_multi_xconnect_ci_master1_result),         //          .result
		.ci_slave_n          (nios2_0_custom_instruction_master_multi_xconnect_ci_master1_n),              //          .n
		.ci_slave_readra     (nios2_0_custom_instruction_master_multi_xconnect_ci_master1_readra),         //          .readra
		.ci_slave_readrb     (nios2_0_custom_instruction_master_multi_xconnect_ci_master1_readrb),         //          .readrb
		.ci_slave_writerc    (nios2_0_custom_instruction_master_multi_xconnect_ci_master1_writerc),        //          .writerc
		.ci_slave_a          (nios2_0_custom_instruction_master_multi_xconnect_ci_master1_a),              //          .a
		.ci_slave_b          (nios2_0_custom_instruction_master_multi_xconnect_ci_master1_b),              //          .b
		.ci_slave_c          (nios2_0_custom_instruction_master_multi_xconnect_ci_master1_c),              //          .c
		.ci_slave_ipending   (nios2_0_custom_instruction_master_multi_xconnect_ci_master1_ipending),       //          .ipending
		.ci_slave_estatus    (nios2_0_custom_instruction_master_multi_xconnect_ci_master1_estatus),        //          .estatus
		.ci_slave_clk        (nios2_0_custom_instruction_master_multi_xconnect_ci_master1_clk),            //          .clk
		.ci_slave_clken      (nios2_0_custom_instruction_master_multi_xconnect_ci_master1_clk_en),         //          .clk_en
		.ci_slave_reset_req  (nios2_0_custom_instruction_master_multi_xconnect_ci_master1_reset_req),      //          .reset_req
		.ci_slave_reset      (nios2_0_custom_instruction_master_multi_xconnect_ci_master1_reset),          //          .reset
		.ci_slave_start      (nios2_0_custom_instruction_master_multi_xconnect_ci_master1_start),          //          .start
		.ci_slave_done       (nios2_0_custom_instruction_master_multi_xconnect_ci_master1_done),           //          .done
		.ci_master_dataa     (nios2_0_custom_instruction_master_multi_slave_translator1_ci_master_dataa),  // ci_master.dataa
		.ci_master_datab     (nios2_0_custom_instruction_master_multi_slave_translator1_ci_master_datab),  //          .datab
		.ci_master_result    (nios2_0_custom_instruction_master_multi_slave_translator1_ci_master_result), //          .result
		.ci_master_n         (nios2_0_custom_instruction_master_multi_slave_translator1_ci_master_n),      //          .n
		.ci_master_clk       (nios2_0_custom_instruction_master_multi_slave_translator1_ci_master_clk),    //          .clk
		.ci_master_clken     (nios2_0_custom_instruction_master_multi_slave_translator1_ci_master_clk_en), //          .clk_en
		.ci_master_reset     (nios2_0_custom_instruction_master_multi_slave_translator1_ci_master_reset),  //          .reset
		.ci_master_start     (nios2_0_custom_instruction_master_multi_slave_translator1_ci_master_start),  //          .start
		.ci_master_done      (nios2_0_custom_instruction_master_multi_slave_translator1_ci_master_done),   //          .done
		.ci_master_readra    (),                                                                           // (terminated)
		.ci_master_readrb    (),                                                                           // (terminated)
		.ci_master_writerc   (),                                                                           // (terminated)
		.ci_master_a         (),                                                                           // (terminated)
		.ci_master_b         (),                                                                           // (terminated)
		.ci_master_c         (),                                                                           // (terminated)
		.ci_master_ipending  (),                                                                           // (terminated)
		.ci_master_estatus   (),                                                                           // (terminated)
		.ci_master_reset_req ()                                                                            // (terminated)
	);

	nios2_mm_interconnect_0 mm_interconnect_0 (
		.pll_0_outclk0_clk                         (pll_0_outclk0_clk),                   //                       pll_0_outclk0.clk
		.arbit_0_reset_reset_bridge_in_reset_reset (rst_controller_reset_out_reset),      // arbit_0_reset_reset_bridge_in_reset.reset
		.arbit_0_avalon_master_address             (arbit_0_avalon_master_address),       //               arbit_0_avalon_master.address
		.arbit_0_avalon_master_waitrequest         (arbit_0_avalon_master_waitrequest),   //                                    .waitrequest
		.arbit_0_avalon_master_chipselect          (arbit_0_avalon_master_chipselect),    //                                    .chipselect
		.arbit_0_avalon_master_read                (arbit_0_avalon_master_read),          //                                    .read
		.arbit_0_avalon_master_readdata            (arbit_0_avalon_master_readdata),      //                                    .readdata
		.arbit_0_avalon_master_write               (arbit_0_avalon_master_write),         //                                    .write
		.arbit_0_avalon_master_writedata           (arbit_0_avalon_master_writedata),     //                                    .writedata
		.mem_s2_address                            (mm_interconnect_0_mem_s2_address),    //                              mem_s2.address
		.mem_s2_write                              (mm_interconnect_0_mem_s2_write),      //                                    .write
		.mem_s2_readdata                           (mm_interconnect_0_mem_s2_readdata),   //                                    .readdata
		.mem_s2_writedata                          (mm_interconnect_0_mem_s2_writedata),  //                                    .writedata
		.mem_s2_byteenable                         (mm_interconnect_0_mem_s2_byteenable), //                                    .byteenable
		.mem_s2_chipselect                         (mm_interconnect_0_mem_s2_chipselect), //                                    .chipselect
		.mem_s2_clken                              (mm_interconnect_0_mem_s2_clken)       //                                    .clken
	);

	nios2_mm_interconnect_1 mm_interconnect_1 (
		.pll_0_outclk0_clk                                 (pll_0_outclk0_clk),                                                   //                       pll_0_outclk0.clk
		.nios2_0_reset_reset_bridge_in_reset_reset         (rst_controller_reset_out_reset),                                      // nios2_0_reset_reset_bridge_in_reset.reset
		.nios2_0_data_master_address                       (nios2_0_data_master_address),                                         //                 nios2_0_data_master.address
		.nios2_0_data_master_waitrequest                   (nios2_0_data_master_waitrequest),                                     //                                    .waitrequest
		.nios2_0_data_master_byteenable                    (nios2_0_data_master_byteenable),                                      //                                    .byteenable
		.nios2_0_data_master_read                          (nios2_0_data_master_read),                                            //                                    .read
		.nios2_0_data_master_readdata                      (nios2_0_data_master_readdata),                                        //                                    .readdata
		.nios2_0_data_master_readdatavalid                 (nios2_0_data_master_readdatavalid),                                   //                                    .readdatavalid
		.nios2_0_data_master_write                         (nios2_0_data_master_write),                                           //                                    .write
		.nios2_0_data_master_writedata                     (nios2_0_data_master_writedata),                                       //                                    .writedata
		.nios2_0_data_master_debugaccess                   (nios2_0_data_master_debugaccess),                                     //                                    .debugaccess
		.nios2_0_instruction_master_address                (nios2_0_instruction_master_address),                                  //          nios2_0_instruction_master.address
		.nios2_0_instruction_master_waitrequest            (nios2_0_instruction_master_waitrequest),                              //                                    .waitrequest
		.nios2_0_instruction_master_read                   (nios2_0_instruction_master_read),                                     //                                    .read
		.nios2_0_instruction_master_readdata               (nios2_0_instruction_master_readdata),                                 //                                    .readdata
		.nios2_0_instruction_master_readdatavalid          (nios2_0_instruction_master_readdatavalid),                            //                                    .readdatavalid
		.jtaguart_0_avalon_jtag_slave_address              (mm_interconnect_1_jtaguart_0_avalon_jtag_slave_address),              //        jtaguart_0_avalon_jtag_slave.address
		.jtaguart_0_avalon_jtag_slave_write                (mm_interconnect_1_jtaguart_0_avalon_jtag_slave_write),                //                                    .write
		.jtaguart_0_avalon_jtag_slave_read                 (mm_interconnect_1_jtaguart_0_avalon_jtag_slave_read),                 //                                    .read
		.jtaguart_0_avalon_jtag_slave_readdata             (mm_interconnect_1_jtaguart_0_avalon_jtag_slave_readdata),             //                                    .readdata
		.jtaguart_0_avalon_jtag_slave_writedata            (mm_interconnect_1_jtaguart_0_avalon_jtag_slave_writedata),            //                                    .writedata
		.jtaguart_0_avalon_jtag_slave_waitrequest          (mm_interconnect_1_jtaguart_0_avalon_jtag_slave_waitrequest),          //                                    .waitrequest
		.jtaguart_0_avalon_jtag_slave_chipselect           (mm_interconnect_1_jtaguart_0_avalon_jtag_slave_chipselect),           //                                    .chipselect
		.mem_s1_address                                    (mm_interconnect_1_mem_s1_address),                                    //                              mem_s1.address
		.mem_s1_write                                      (mm_interconnect_1_mem_s1_write),                                      //                                    .write
		.mem_s1_readdata                                   (mm_interconnect_1_mem_s1_readdata),                                   //                                    .readdata
		.mem_s1_writedata                                  (mm_interconnect_1_mem_s1_writedata),                                  //                                    .writedata
		.mem_s1_byteenable                                 (mm_interconnect_1_mem_s1_byteenable),                                 //                                    .byteenable
		.mem_s1_chipselect                                 (mm_interconnect_1_mem_s1_chipselect),                                 //                                    .chipselect
		.mem_s1_clken                                      (mm_interconnect_1_mem_s1_clken),                                      //                                    .clken
		.nios2_0_debug_mem_slave_address                   (mm_interconnect_1_nios2_0_debug_mem_slave_address),                   //             nios2_0_debug_mem_slave.address
		.nios2_0_debug_mem_slave_write                     (mm_interconnect_1_nios2_0_debug_mem_slave_write),                     //                                    .write
		.nios2_0_debug_mem_slave_read                      (mm_interconnect_1_nios2_0_debug_mem_slave_read),                      //                                    .read
		.nios2_0_debug_mem_slave_readdata                  (mm_interconnect_1_nios2_0_debug_mem_slave_readdata),                  //                                    .readdata
		.nios2_0_debug_mem_slave_writedata                 (mm_interconnect_1_nios2_0_debug_mem_slave_writedata),                 //                                    .writedata
		.nios2_0_debug_mem_slave_byteenable                (mm_interconnect_1_nios2_0_debug_mem_slave_byteenable),                //                                    .byteenable
		.nios2_0_debug_mem_slave_waitrequest               (mm_interconnect_1_nios2_0_debug_mem_slave_waitrequest),               //                                    .waitrequest
		.nios2_0_debug_mem_slave_debugaccess               (mm_interconnect_1_nios2_0_debug_mem_slave_debugaccess),               //                                    .debugaccess
		.performance_counter_0_control_slave_address       (mm_interconnect_1_performance_counter_0_control_slave_address),       // performance_counter_0_control_slave.address
		.performance_counter_0_control_slave_write         (mm_interconnect_1_performance_counter_0_control_slave_write),         //                                    .write
		.performance_counter_0_control_slave_readdata      (mm_interconnect_1_performance_counter_0_control_slave_readdata),      //                                    .readdata
		.performance_counter_0_control_slave_writedata     (mm_interconnect_1_performance_counter_0_control_slave_writedata),     //                                    .writedata
		.performance_counter_0_control_slave_begintransfer (mm_interconnect_1_performance_counter_0_control_slave_begintransfer), //                                    .begintransfer
		.sys_clk_timer_s1_address                          (mm_interconnect_1_sys_clk_timer_s1_address),                          //                    sys_clk_timer_s1.address
		.sys_clk_timer_s1_write                            (mm_interconnect_1_sys_clk_timer_s1_write),                            //                                    .write
		.sys_clk_timer_s1_readdata                         (mm_interconnect_1_sys_clk_timer_s1_readdata),                         //                                    .readdata
		.sys_clk_timer_s1_writedata                        (mm_interconnect_1_sys_clk_timer_s1_writedata),                        //                                    .writedata
		.sys_clk_timer_s1_chipselect                       (mm_interconnect_1_sys_clk_timer_s1_chipselect),                       //                                    .chipselect
		.sysid_control_slave_address                       (mm_interconnect_1_sysid_control_slave_address),                       //                 sysid_control_slave.address
		.sysid_control_slave_readdata                      (mm_interconnect_1_sysid_control_slave_readdata)                       //                                    .readdata
	);

	nios2_irq_mapper irq_mapper (
		.clk           (pll_0_outclk0_clk),              //       clk.clk
		.reset         (rst_controller_reset_out_reset), // clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq),       // receiver0.irq
		.receiver1_irq (irq_mapper_receiver1_irq),       // receiver1.irq
		.sender_irq    (nios2_0_irq_irq)                 //    sender.irq
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~reset_reset_n),                     // reset_in0.reset
		.clk            (pll_0_outclk0_clk),                  //       clk.clk
		.reset_out      (rst_controller_reset_out_reset),     // reset_out.reset
		.reset_req      (rst_controller_reset_out_reset_req), //          .reset_req
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_in1      (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

endmodule
